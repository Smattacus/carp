`define NUM_TEST_VECS 1


package clock; 
    parameter time period = 8ns;
endpackage : clock
